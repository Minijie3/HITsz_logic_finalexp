`timescale 1ns / 1ps

module led_list(
    input [7:0] num,
    output reg [7:0] SEGS
);
    always @* begin
        case(num)
            48: SEGS <= 8'b00000011; //00110000：0
            49: SEGS <= 8'b10011111; //00110001：1
            50: SEGS <= 8'b00100101; //00110010：2
            51: SEGS <= 8'b00001101; //00110011：3
            52: SEGS <= 8'b10011001; //00110100：4
            53: SEGS <= 8'b01001001; //00110101：5
            54: SEGS <= 8'b01000001; //00110110：6
            55: SEGS <= 8'b00011111; //00110111：7
            56: SEGS <= 8'b00000001; //00111000：8
            57: SEGS <= 8'b00001001; //00111001：9
            65: SEGS <= 8'b00010001; //01000001：A
            66: SEGS <= 8'b11000001; //01000010：B
            67: SEGS <= 8'b11100101; //01000011：C
            68: SEGS <= 8'b10000101; //01000100：D
            69: SEGS <= 8'b01100001; //01000101：E
            70: SEGS <= 8'b01110001; //01000110：F
            default: SEGS <= 8'b11111111; //0-F 之外的统一不显示
        endcase
    end
endmodule